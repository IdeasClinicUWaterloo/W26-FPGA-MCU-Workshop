library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY activity_2 IS
    PORT (
        SW : IN STD_LOGIC_VECTOR(3 DOWNTO 0);    -- SWITCH DECLARATION
        HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)	 -- SEVEN SEGMENT OUTPUT
    );
END activity_2;

ARCHITECTURE Behavioral OF activity_2 IS
   
	-- SIGNAL declaration

	
    
BEGIN

    --PROCESS declaration
	 
	 
	 


	 --PROCESS end
    
	 --HEX0 assignment

	 
    
END Behavioral;