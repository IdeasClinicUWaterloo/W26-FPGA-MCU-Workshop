-- ========================================
-- ACTIVITY 3: activity_3.vhd
-- Full Adder with Seven-Segment Display
-- ========================================
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity activity_3 is
   Port (
       SW : in STD_LOGIC_VECTOR(2 downto 0);    -- SW0=A, SW1=B, SW2=Cin
       HEX1 : out STD_LOGIC_VECTOR(6 downto 0)
   );
end activity_3;

architecture Behavioral of activity_3 is
    
	--SIGNAL declarations

    
begin
    
   -- Full Adder Logic

	
   
	
	-- Convert Full Adder Result to 7-segment display
    
	 
	 
	 
	-- HEX1 assignment
	 
    
end Behavioral;