-- ========================================
-- ACTIVITY 1: activity_1.vhd
-- Full Adder - outputs to LEDs
-- ========================================
library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY activity_1 IS
    PORT (
        SW : IN STD_LOGIC_VECTOR(2 downto 0);   -- SW(0) = A, SW(1) = B, SW(2) = C
        LED : OUT STD_LOGIC_VECTOR(1 downto 0)  -- LED(0) = SUM, LED(1) = CARRY
    );
END activity_1;

architecture Behavioral of activity_1 is
	
	--SIGNAL declarations
	
	

BEGIN
	

	
	
	-- LED assignments

	
	 
END Behavioral;